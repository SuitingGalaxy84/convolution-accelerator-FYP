`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: University of Electronic Science and Technology of China
// Engineer: Sun Yucheng
// 
// Create Date: XX
// Design Name: PE Key-Lock Checker 
// Module Name: SV_DummyPE_KL
// Project Name: A Convolution Accelerator for PyTorch Deep Learning Framework
// Target Devices: PYNQ Z1
// Tool Versions: Vivado 20XX.XX
// Description: 
/*
    a LOCK-KEY scheme is created. Every PE is assgined with a unique ROW-COL tag at the initialization. The PE
    can be activated only when the corresponding ROW-COL tag is provided. This facilitates an efficient control
    of the PE array.
 */
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////
`include "interface.sv"

module caster#(
    parameter DATA_WIDTH = 16,
    parameter NUM_COL = 4
)(
    input wire clk,
    input wire rstn,

    CASTER_IF.CASTER_data CASTER_data,
    CASTER_IF.CASTER_ctrl CASTER_ctrl
    );

    reg [$clog2(NUM_COL)-1:0] caster_id; 
    always_ff @(posedge clk or negedge rstn) begin // facilitate the PE matching
        if(~rstn) begin
            caster_id <= 0;
        end else begin
            caster_id <= CASTER_ctrl.ID;
        end 
    end

    always_comb begin: PE_to_BUS//facilitate hte data output from PE to bus
        case ({CASTER_ctrl.PE_VALID, CASTER_ctrl.CASTER_EN, (CASTER_ctrl.TAG == caster_id ? 1'b1 : 1'b0)})
            3'b111 : begin 
                CASTER_data.data_C2B = CASTER_data.data_C2P;
            end 
            default: begin 
                CASTER_data.data_C2B = 0;
            end 
        endcase
        CASTER_ctrl.CASTER_VALID = CASTER_ctrl.PE_VALID; // notify the BUS that the PE has valid data
    end

    always_comb begin : BUS_to_PE//facilitate the data input from bus to PE
        case ({CASTER_ctrl.PE_READY, CASTER_ctrl.CASTER_EN, (CASTER_ctrl.TAG == caster_id ? 1'b1 : 1'b0)})
            3'b111 : begin 
                CASTER_ctrl.PE_EN = 1'b1;
                CASTER_data.data_C2P = CASTER_data.data_B2C;
            end 
            default: begin 
                CASTER_ctrl.PE_EN = 1'b0;
                CASTER_data.data_C2P = 0;
            end
        endcase
        CASTER_ctrl.CASTER_READY = CASTER_ctrl.PE_READY; // notify the BUS that the PE is ready to accept data
    end







endmodule