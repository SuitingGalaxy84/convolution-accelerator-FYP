`include "def.sv"


module SV_PE_link #(
    parameter DATA_WIDTH = 16,
    parameter NUM_ROW = 3,
    parameter NUM_COL = 4
)(

)
    

endmodule