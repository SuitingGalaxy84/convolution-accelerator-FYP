//TODO: design a benchmark for the PE set